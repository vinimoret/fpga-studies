module leds (
    output wire D1,
    output wire D2,
    output wire D3,
    output wire D4,
    output wire D5,
    output wire D6,
    output wire D7,
    output wire D8
);

assign D1 = 1'b0; // Set D1 to high
assign D2 = 1'b0; // Set D2 to low
assign D3 = 1'b0; // Set D2 to low
assign D4 = 1'b0; // Set D2 to low
assign D5 = 1'b0; // Set D2 to low
assign D6 = 1'b0; // Set D2 to low
assign D7 = 1'b0; // Set D2 to low
assign D8 = 1'b0; // Set D2 to low

endmodule